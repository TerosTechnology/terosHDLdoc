package mynewpackage is
    
end package;