process (all)
begin
    
end process;