library ieee;
use ieee.std_logic_1164.all;

package mytypes is
    type main_sm_type is (IDLE,PUSHA,PUSHB,FINISH); --! main state machine states 
end package;