module tb_mytb(
    input clk,
    input rstn
);

mymodule dut(
    .rstn (rstn),
    .clk (clk)
);


endmodule
