module myconsts ();

localparam SN=11223344; //! SN for this node
    
endmodule