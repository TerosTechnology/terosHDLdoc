entity ports is
    port (
        clk   : in std_logic; --! my clock
        reset : in std_logic --! reset of everything
    );
end entity;