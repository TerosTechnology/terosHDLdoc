library ieee;
use ieee.std_logic_1164.all;
package mypackage is
    function func1 (x:integer) return std_logic;
    
end package;
package body mypackage is
    function func1 (x:integer) return std_logic is
    begin
        
    end function;
end package body;