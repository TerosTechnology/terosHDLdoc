module funcs ;

function reg[1:0] myfunc(input a,b);

    myfunc = {a,b};
endfunction


endmodule

