--! Entity example
-- description
entity entity is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity;