library ieee;
use ieee.std_logic_1164.all;

package mytypes is
    type t_my_custom_type is range 0 to 1000; --! my custom type description
end package;