//! AXI-4 Stream
typedef struct packed {  
    logic [7:0] data;
    logic [0:0] valid;
    logic [0:0] clk;
} mystruct;
    
