package mypackage is
    constant DATA_WIDTH : integer := 35; --! number of bits
    constant ADDR_WIDTH : integer := 21; --! number of bits
    
end package;