entity entity is
    port (
        --! Port description 0
        clk   : in std_logic;
        reset : in std_logic --! Port description 1
    );
end entity;